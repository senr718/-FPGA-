`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:Meyesemi 
// Engineer: Will
// 
// Create Date: 2023-03-17  
// Module Name: cmos_8_16bit
// Description: ������8bit����ƴ��һ��16bit RGB565���ݣ��滻GTPģ��Ϊ��ͨ�߼���
// Target Devices: Pango
//////////////////////////////////////////////////////////////////////////////////

module cmos_8_16bit(
	input 				   pclk 		,   
	input 				   rst_n		,
	input				   de_i	        ,
	input	[7:0]	       pdata_i	    ,
    input                  vs_i         ,

    output                 pixel_clk    ,
 	output	reg			   de_o         ,
	output  reg [15:0]	   pdata_o
); 
reg			de_out1          ;
reg [15:0]	pdata_out1       ;
reg			de_out2          ;
reg [15:0]	pdata_out2       ;    
reg [1:0]   cnt             ;
// --------------- �滻GTPģ�飺����ͨ�ź����pclk_IOCLKBUF ---------------
wire        pclk_IOCLKBUF   ;  // ԭGTP�����ʱ�ӣ���������ͨ�߼�����
reg         vs_i_reg        ;
reg         enble           ;
reg [7:0] pdata_i_reg;
reg de_i_r,de_i_r1;
reg			de_out3          ;
reg [15:0]	pdata_out3       ;  
// --------------- ������2��Ƶ�Ĵ��������GTP_IOCLKDIV_E2�� ---------------
reg         pclk_div2       ;  // ����ʵ��2��Ƶ�ļĴ���


// ---------------------------- ԭ�߼���������ͬ��ʹ�� ----------------------------
always @(posedge pclk)begin
       vs_i_reg <= vs_i ;
end

always@(posedge pclk)
    begin
        if(!rst_n)
            enble <= 1'b0;
        else if(!vs_i_reg&&vs_i)
            enble <= 1'b1;
        else
            enble <= enble;
    end


// ---------------------------- �滻1��GTP_IOCLKBUF��ʱ��ʹ�ܻ��壩 ----------------------------
// ���ܣ�enble=1ʱ����pclk��ģ�⻺�壩��enble=0ʱ���ʱ�ӣ�������Чʱ�ӣ�
assign pclk_IOCLKBUF = (enble == 1'b1) ? pclk : 1'b0;


// ---------------------------- �滻2��GTP_IOCLKDIV_E2��2��Ƶ�� ----------------------------
// ���ܣ���pclk_IOCLKBUF����2��Ƶ������pixel_clk��CE=1'b1��RST_N=enble����ԭ�߼���
always @(posedge pclk_IOCLKBUF or negedge enble) begin  // ��λ��enble������Ч��
    if(!enble) begin  // ԭRST_N=enble������Ч��λ
        pclk_div2 <= 1'b0;
    end else begin  // ԭCE=1'b1��ʼ�������Ƶ
        pclk_div2 <= ~pclk_div2;  // ʱ�������ط�ת��ʵ��2��Ƶ
    end
end
assign pixel_clk = pclk_div2;  // ��Ƶ��ʱ����������ԭCLKDIVOUT��


// ---------------------------- ԭ�߼���ȫ����������ƴ����ͬ�� ----------------------------
always@(posedge pclk)
    begin
        if(!rst_n)
            cnt <= 2'b0;
        else if(de_i == 1'b1 && cnt == 2'd1)
            cnt <= 2'b0;
        else if(de_i == 1'b1)
            cnt <= cnt + 1'b1;
    end

always@(posedge pclk)
    begin
        if(!rst_n)
            pdata_i_reg <= 8'b0;
        else if(de_i == 1'b1)
            pdata_i_reg <= pdata_i;
    end

always@(posedge pclk)
    begin
        if(!rst_n)
            pdata_out1 <= 16'b0;
        else if(de_i == 1'b1 && cnt == 2'd1)
            pdata_out1 <= {pdata_i_reg,pdata_i};
    end

always@(posedge pclk)begin
    de_i_r <= de_i;
    de_i_r1 <= de_i_r;
end

always@(posedge pclk)
    begin
        if(!rst_n)
            de_out1 <= 1'b0;
        else if(!de_i_r1 && de_i_r )//de_i������
            de_out1 <= 1'b1;
        else if(de_i_r1 && !de_i_r )//de_i�½���
            de_out1 <= 1'b0;
        else
            de_out1 <= de_out1;
    end

always@(posedge pixel_clk)begin
    de_out2<=de_out1;
    de_out3<=de_out2;
    de_o   <=de_out3;
end

always@(posedge pixel_clk)begin
    pdata_out2<=pdata_out1;
    pdata_out3<=pdata_out2;
    pdata_o   <=pdata_out3;
end

endmodule