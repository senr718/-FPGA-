module fifo_32to128 (
    input               clk_100m,        // ��ʱ��
    input               rst_n,           // ȫ�ָ�λ������Ч��
    input        [31:0] fifo_rd_data,    // FIFO�����32bit����
    input               fifo_empty,      // FIFO�ձ�־���͵�ƽ�ǿգ�
    input               blk_state_WRITE, // �ⲿWRITE״̬������Ч��
    output reg          fifo_rd_en,      // FIFO��ʹ��
    output reg  [127:0] data_128bit,     // ƴ�Ӻ��128bit����
    output reg          data_128_valid   // 128bit������Ч��־
);

reg [1:0] cnt_read;                     // ��ȡ��������0~3����FIFO��ʱ���ֵ�ǰֵ
reg [1:0] next_cnt_read;  
reg [31:0] data_reg [3:0];              // �����ݴ�Ĵ�����FIFO��ʱ��������
localparam IDLE  = 1'b0, READ = 1'b1;
reg current_state, next_state;

// ״̬����ת�����ڡ�����4�����ݡ����˳�WRITE״̬��ʱ����IDLE��FIFO��ʱ����READ
always @(posedge clk_100m or negedge rst_n) begin
    if (!rst_n) current_state <= IDLE;
    else current_state <= next_state;
end

// ״̬����̬�߼���FIFO��ʱ���˳�READ������ͣ��ȡ
always @(*) begin
    case (current_state)
        IDLE: begin
            // ����WRITE״̬��FIFO�ǿ�ʱ������READ
            next_state = (blk_state_WRITE && !fifo_empty) ? READ : IDLE;
        end
        READ: begin
            // �˳�READ��Ψһ����������4������ �� �˳�WRITE״̬����FIFO���޹أ�
            next_state = (cnt_read == 2'd3 || !blk_state_WRITE) ? IDLE : READ;
        end
        default: next_state = IDLE;
    endcase
end

// ��ʹ�ܣ�����READ״̬��FIFO�ǿա�WRITE״̬ʱ��Ч��FIFO��ʱ�Զ�Ϊ0����ͣ��ȡ��
always @(posedge clk_100m or negedge rst_n) begin
    if (!rst_n) fifo_rd_en <= 1'b0;
    else begin
        fifo_rd_en <= (current_state == READ) && !fifo_empty && blk_state_WRITE;
    end
end

// ��������������Ч��ʱ������FIFO��ʱ���ֵ�ǰֵ���˳�WRITEʱ����
always @(posedge clk_100m or negedge rst_n) begin
    if (!rst_n) begin
        cnt_read <= 2'd0;
        next_cnt_read <= 2'd0;
    end else if (!blk_state_WRITE) begin  // �˳�WRITE״̬��ǿ�����㣨������ֹ��
        cnt_read <= 2'd0;
        next_cnt_read <= 2'd0;
    end else if (fifo_rd_en) begin  // ��Ч��ʱ����������FIFO�ǿ�����READ״̬��
        cnt_read <= next_cnt_read + 2'd1;
        next_cnt_read <= next_cnt_read + 2'd1;
    end
    // �����߼���FIFO��ʱ��fifo_rd_en=0����cnt_read���ֵ�ǰֵ�������㣩
end

// ���ݼĴ�����FIFO��ʱ�������ݣ���Ч��ʱ�洢���˳�WRITEʱ����
always @(posedge clk_100m or negedge rst_n) begin
    if (!rst_n) begin
        data_reg[0] <= 32'd0;
        data_reg[1] <= 32'd0;
        data_reg[2] <= 32'd0;
        data_reg[3] <= 32'd0;
    end else if (!blk_state_WRITE) begin  // �˳�WRITE״̬���������ݣ�������ֹ��
        data_reg[0] <= 32'd0;
        data_reg[1] <= 32'd0;
        data_reg[2] <= 32'd0;
        data_reg[3] <= 32'd0;
    end else if (fifo_rd_en) begin  // ��Ч��ʱ�洢���ݣ�FIFO�ǿ�ʱ������䣩
        case (cnt_read)
            2'd0: data_reg[0] <= fifo_rd_data;
            2'd1: data_reg[1] <= fifo_rd_data;
            2'd2: data_reg[2] <= fifo_rd_data;
            2'd3: data_reg[3] <= fifo_rd_data;
        endcase
    end
    // �����߼���FIFO��ʱ��data_reg�����Ѵ����ݣ��������
end

// 128bit������Ч������4������ȫ������ʱ��Ч
always @(posedge clk_100m or negedge rst_n) begin
    if (!rst_n) begin
        data_128bit <= 128'd0;
        data_128_valid <= 1'b0;
    end else begin
        // �������4�����ݣ�cnt_read=3�Ҷ�ʹ����Ч�������128bit����
        if (cnt_read == 2'd3 && fifo_rd_en) begin
            data_128bit <= {data_reg[3], data_reg[2], data_reg[1], data_reg[0]};
            data_128_valid <= 1'b1;
        end else begin
            data_128_valid <= 1'b0;
        end
    end
end

endmodule