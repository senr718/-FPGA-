//���Լ򵥵����ݽ���
//����i2cSlave_define.v���޸�IIC��ַ
//��registerInterface.v���޸ļĴ���
module iic_slave_top
(
    input    wire            sys_clk    ,   //ϵͳʱ�� 25MHZ

	input	 wire		     i2c_scl    ,	// IIC ʱ����
	inout 	 wire		     i2c_sda    ,	// IIC ������
	output	 wire    [1:0]	 led            // �û�LED

);
//IIC register                                   
wire  [7:0]led_reg;//0x01
wire  [7:0] myReg0_flag;

wire    clk_100m    ;
wire    rst_n       ;
reg   Reg0_wr_en;
reg   Reg1_wr_en;
reg   [7:0]  myReg0_w;
reg   [7:0]  myReg1_w;
//����100MHZ��ʱ��
iic_pll iic_pll_inst (
  .clkout0(clk_100m),    // output
  .lock(rst_n),          // output
  .clkin1(sys_clk)       // input
);
//iic slaveģ��
i2cSlave i2cSlave_u (
	.clk		(clk_100m),		
	.rst		(~rst_n  ),		
	.sda		(i2c_sda ),		
	.scl		(i2c_scl ),	
    .Reg0_wr_en (Reg0_wr_en ),		
    .Reg1_wr_en (Reg1_wr_en ),		
    .myReg0_w   (myReg0_w ),		
	.myReg1_w   (myReg1_w ),		
	.myReg0		(myReg0_flag ),		
	.myReg1		(led_reg )		
);
//����01�Ĵ����ĵ�2bit
assign	led 	= led_reg[1:0];




endmodule