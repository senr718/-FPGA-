module rgb565_to_rgb888 (
    input                  rst_n,       // ���븴λ������߼��½����ڸ�λʱ���㣩
    input        [15:0]    i_rgb565,    // ����RGB565����
    output       [23:0]    o_rgb888    // ���RGB888���ݣ�R[23:16],G[15:8],B[7:0]��

);

// ����߼�ʵ�֣���ʱ���ӳ٣����������ͬ���仯
assign o_rgb888 = (!rst_n) ? 24'd0 : 
                 {i_rgb565[15:11], 3'b000,  // R: 5bit��8bit����3��0��
                  i_rgb565[10:5],  2'b00,   // G: 6bit��8bit����2��0��
                  i_rgb565[4:0],   3'b000}; // B: 5bit��8bit����3��0��

endmodule